module xor_mod (A,B,Y);
    output Y;
    input A,B;

    xor(Y,A,B);
endmodule